// Code your testbench here
// or browse Examples
`include "eth_testbench_top.sv"