interface mux_intf();
	logic x;
	logic y;
  	logic v;
	logic z;
    logic [1:0]select;
	logic mux_out;
endinterface
