interface intf();
  
  //declaring the signals
  logic [3:0] a;
  logic [3:0] b;
  logic [7:0] c;
  
 
 // modport driver (output a, b, input c);
  
endinterface