interface intf();
  
  //declaring the signals
  logic [3:0] a;
  logic [3:0] b;
  logic sel;
  logic [3:0] out;
  
  
 
  
endinterface