class generator;
  rand transaction trans;
  
  
  mailbox gen2driv;
  
  
  function new(mailbox gen2driv);
    this.gen2driv = gen2driv;
  endfunction
  
  task run;
      trans=new();
    begin
      trans.constraint_mode(0);
      trans.c_Y8.constraint_mode(1); 
      if( !trans.randomize()) 
        $error("Gen::trans randomization failed");
      //assert(trans.randomize());
      trans.display("[ Generator ] ");
      gen2driv.put(trans);
    end
  endtask
  
endclass:generator
      
      
    
  