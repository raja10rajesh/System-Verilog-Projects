interface mux_intf();
	logic x;
	logic y;
	logic select;
	logic mux_out;
endinterface
