interface intf();
  
  //declaring the signals
  logic [2:0] in;
  logic [7:0] out;
  logic en;
  

  
endinterface