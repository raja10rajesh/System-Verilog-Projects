// Code your design here
`include "simpleadder.v"