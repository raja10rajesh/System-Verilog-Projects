interface intf();
  
  //declaring the signals
  logic [7:0] Y;
  logic [2:0] out;

  

  
endinterface